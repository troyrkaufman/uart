// fifo.sv
// Troy Kaufman
// 